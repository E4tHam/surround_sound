
/* delaydampener.v */


module Dampener (
    input     [7:0] theta       ,
    output    [7:0] damp
);

    assign damp  = 0;

endmodule
